// sopc.v

// Generated using ACDS version 13.1 162 at 2018.11.20.16:59:48

`timescale 1 ps / 1 ps
module sopc (
		input  wire        reset_n,                   //             clk_clk_in_reset.reset_n
		output wire        out_port_from_the_LAN_RST, //  LAN_RST_external_connection.export
		output wire        out_port_from_the_LAN_CS,  //   LAN_CS_external_connection.export
		input  wire        MISO_to_the_LAN,           //                 LAN_external.MISO
		output wire        MOSI_from_the_LAN,         //                             .MOSI
		output wire        SCLK_from_the_LAN,         //                             .SCLK
		output wire        SS_n_from_the_LAN,         //                             .SS_n
		input  wire        clk,                       //                   clk_clk_in.clk
		input  wire        in_port_to_the_LAN_NINT,   // LAN_NINT_external_connection.export
		output wire        dclk_from_the_epcs,        //                epcs_external.dclk
		output wire        sce_from_the_epcs,         //                             .sce
		output wire        sdo_from_the_epcs,         //                             .sdo
		input  wire        data0_to_the_epcs,         //                             .data0
		input  wire [31:0] time_export,               //                         time.export
		input  wire [31:0] ch1_count_export,          //                    ch1_count.export
		output wire [7:0]  addr_export,               //                         addr.export
		input  wire [7:0]  rdata_export,              //                        rdata.export
		output wire [7:0]  wdata_export,              //                        wdata.export
		output wire [7:0]  signals_export,            //                      signals.export
		input  wire [7:0]  status_export,             //                       status.export
		output wire [31:0] wdata32_export,            //                      wdata32.export
		output wire [31:0] rdata32_export,            //                      rdata32.export
		input  wire [31:0] ch2_count_export,          //                    ch2_count.export
		input  wire [31:0] ch3_count_export,          //                    ch3_count.export
		input  wire [31:0] ch4_count_export           //                    ch4_count.export
	);

	wire  [31:0] mm_interconnect_0_onchip_mem_s1_writedata;                 // mm_interconnect_0:onchip_mem_s1_writedata -> onchip_mem:writedata
	wire  [13:0] mm_interconnect_0_onchip_mem_s1_address;                   // mm_interconnect_0:onchip_mem_s1_address -> onchip_mem:address
	wire         mm_interconnect_0_onchip_mem_s1_chipselect;                // mm_interconnect_0:onchip_mem_s1_chipselect -> onchip_mem:chipselect
	wire         mm_interconnect_0_onchip_mem_s1_clken;                     // mm_interconnect_0:onchip_mem_s1_clken -> onchip_mem:clken
	wire         mm_interconnect_0_onchip_mem_s1_write;                     // mm_interconnect_0:onchip_mem_s1_write -> onchip_mem:write
	wire  [31:0] mm_interconnect_0_onchip_mem_s1_readdata;                  // onchip_mem:readdata -> mm_interconnect_0:onchip_mem_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_mem_s1_byteenable;                // mm_interconnect_0:onchip_mem_s1_byteenable -> onchip_mem:byteenable
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [17:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire   [1:0] mm_interconnect_0_pio_count3_s1_address;                   // mm_interconnect_0:pio_count3_s1_address -> pio_count3:address
	wire  [31:0] mm_interconnect_0_pio_count3_s1_readdata;                  // pio_count3:readdata -> mm_interconnect_0:pio_count3_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_time_s1_address;                     // mm_interconnect_0:pio_time_s1_address -> pio_time:address
	wire  [31:0] mm_interconnect_0_pio_time_s1_readdata;                    // pio_time:readdata -> mm_interconnect_0:pio_time_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_signals_0_s1_address;                // mm_interconnect_0:pio_signals_0_s1_address -> pio_signals_0:address
	wire  [31:0] mm_interconnect_0_pio_signals_0_s1_readdata;               // pio_signals_0:readdata -> mm_interconnect_0:pio_signals_0_s1_readdata
	wire  [15:0] mm_interconnect_0_lan_spi_control_port_writedata;          // mm_interconnect_0:LAN_spi_control_port_writedata -> LAN:data_from_cpu
	wire   [2:0] mm_interconnect_0_lan_spi_control_port_address;            // mm_interconnect_0:LAN_spi_control_port_address -> LAN:mem_addr
	wire         mm_interconnect_0_lan_spi_control_port_chipselect;         // mm_interconnect_0:LAN_spi_control_port_chipselect -> LAN:spi_select
	wire         mm_interconnect_0_lan_spi_control_port_write;              // mm_interconnect_0:LAN_spi_control_port_write -> LAN:write_n
	wire         mm_interconnect_0_lan_spi_control_port_read;               // mm_interconnect_0:LAN_spi_control_port_read -> LAN:read_n
	wire  [15:0] mm_interconnect_0_lan_spi_control_port_readdata;           // LAN:data_to_cpu -> mm_interconnect_0:LAN_spi_control_port_readdata
	wire   [1:0] mm_interconnect_0_pio_count4_s1_address;                   // mm_interconnect_0:pio_count4_s1_address -> pio_count4:address
	wire  [31:0] mm_interconnect_0_pio_count4_s1_readdata;                  // pio_count4:readdata -> mm_interconnect_0:pio_count4_s1_readdata
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_writedata;        // mm_interconnect_0:epcs_epcs_control_port_writedata -> epcs:writedata
	wire   [8:0] mm_interconnect_0_epcs_epcs_control_port_address;          // mm_interconnect_0:epcs_epcs_control_port_address -> epcs:address
	wire         mm_interconnect_0_epcs_epcs_control_port_chipselect;       // mm_interconnect_0:epcs_epcs_control_port_chipselect -> epcs:chipselect
	wire         mm_interconnect_0_epcs_epcs_control_port_write;            // mm_interconnect_0:epcs_epcs_control_port_write -> epcs:write_n
	wire         mm_interconnect_0_epcs_epcs_control_port_read;             // mm_interconnect_0:epcs_epcs_control_port_read -> epcs:read_n
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_readdata;         // epcs:readdata -> mm_interconnect_0:epcs_epcs_control_port_readdata
	wire   [1:0] mm_interconnect_0_pio_count2_s1_address;                   // mm_interconnect_0:pio_count2_s1_address -> pio_count2:address
	wire  [31:0] mm_interconnect_0_pio_count2_s1_readdata;                  // pio_count2:readdata -> mm_interconnect_0:pio_count2_s1_readdata
	wire  [31:0] mm_interconnect_0_data32_in_s1_writedata;                  // mm_interconnect_0:data32_in_s1_writedata -> data32_in:writedata
	wire   [1:0] mm_interconnect_0_data32_in_s1_address;                    // mm_interconnect_0:data32_in_s1_address -> data32_in:address
	wire         mm_interconnect_0_data32_in_s1_chipselect;                 // mm_interconnect_0:data32_in_s1_chipselect -> data32_in:chipselect
	wire         mm_interconnect_0_data32_in_s1_write;                      // mm_interconnect_0:data32_in_s1_write -> data32_in:write_n
	wire  [31:0] mm_interconnect_0_data32_in_s1_readdata;                   // data32_in:readdata -> mm_interconnect_0:data32_in_s1_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [17:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                               // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire  [31:0] mm_interconnect_0_pio_addr_s1_writedata;                   // mm_interconnect_0:pio_addr_s1_writedata -> pio_addr:writedata
	wire   [1:0] mm_interconnect_0_pio_addr_s1_address;                     // mm_interconnect_0:pio_addr_s1_address -> pio_addr:address
	wire         mm_interconnect_0_pio_addr_s1_chipselect;                  // mm_interconnect_0:pio_addr_s1_chipselect -> pio_addr:chipselect
	wire         mm_interconnect_0_pio_addr_s1_write;                       // mm_interconnect_0:pio_addr_s1_write -> pio_addr:write_n
	wire  [31:0] mm_interconnect_0_pio_addr_s1_readdata;                    // pio_addr:readdata -> mm_interconnect_0:pio_addr_s1_readdata
	wire   [1:0] mm_interconnect_0_lan_nint_s1_address;                     // mm_interconnect_0:LAN_NINT_s1_address -> LAN_NINT:address
	wire  [31:0] mm_interconnect_0_lan_nint_s1_readdata;                    // LAN_NINT:readdata -> mm_interconnect_0:LAN_NINT_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_wdata_s1_writedata;                  // mm_interconnect_0:pio_wdata_s1_writedata -> pio_wdata:writedata
	wire   [1:0] mm_interconnect_0_pio_wdata_s1_address;                    // mm_interconnect_0:pio_wdata_s1_address -> pio_wdata:address
	wire         mm_interconnect_0_pio_wdata_s1_chipselect;                 // mm_interconnect_0:pio_wdata_s1_chipselect -> pio_wdata:chipselect
	wire         mm_interconnect_0_pio_wdata_s1_write;                      // mm_interconnect_0:pio_wdata_s1_write -> pio_wdata:write_n
	wire  [31:0] mm_interconnect_0_pio_wdata_s1_readdata;                   // pio_wdata:readdata -> mm_interconnect_0:pio_wdata_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_count_s1_address;                    // mm_interconnect_0:pio_count_s1_address -> pio_count:address
	wire  [31:0] mm_interconnect_0_pio_count_s1_readdata;                   // pio_count:readdata -> mm_interconnect_0:pio_count_s1_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;       // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;           // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;             // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;              // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;          // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_data32_s1_writedata;                     // mm_interconnect_0:data32_s1_writedata -> data32:writedata
	wire   [1:0] mm_interconnect_0_data32_s1_address;                       // mm_interconnect_0:data32_s1_address -> data32:address
	wire         mm_interconnect_0_data32_s1_chipselect;                    // mm_interconnect_0:data32_s1_chipselect -> data32:chipselect
	wire         mm_interconnect_0_data32_s1_write;                         // mm_interconnect_0:data32_s1_write -> data32:write_n
	wire  [31:0] mm_interconnect_0_data32_s1_readdata;                      // data32:readdata -> mm_interconnect_0:data32_s1_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [1:0] mm_interconnect_0_pio_rdata_s1_address;                    // mm_interconnect_0:pio_rdata_s1_address -> pio_rdata:address
	wire  [31:0] mm_interconnect_0_pio_rdata_s1_readdata;                   // pio_rdata:readdata -> mm_interconnect_0:pio_rdata_s1_readdata
	wire  [31:0] mm_interconnect_0_lan_cs_s1_writedata;                     // mm_interconnect_0:LAN_CS_s1_writedata -> LAN_CS:writedata
	wire   [1:0] mm_interconnect_0_lan_cs_s1_address;                       // mm_interconnect_0:LAN_CS_s1_address -> LAN_CS:address
	wire         mm_interconnect_0_lan_cs_s1_chipselect;                    // mm_interconnect_0:LAN_CS_s1_chipselect -> LAN_CS:chipselect
	wire         mm_interconnect_0_lan_cs_s1_write;                         // mm_interconnect_0:LAN_CS_s1_write -> LAN_CS:write_n
	wire  [31:0] mm_interconnect_0_lan_cs_s1_readdata;                      // LAN_CS:readdata -> mm_interconnect_0:LAN_CS_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_signals_s1_writedata;                // mm_interconnect_0:pio_signals_s1_writedata -> pio_signals:writedata
	wire   [1:0] mm_interconnect_0_pio_signals_s1_address;                  // mm_interconnect_0:pio_signals_s1_address -> pio_signals:address
	wire         mm_interconnect_0_pio_signals_s1_chipselect;               // mm_interconnect_0:pio_signals_s1_chipselect -> pio_signals:chipselect
	wire         mm_interconnect_0_pio_signals_s1_write;                    // mm_interconnect_0:pio_signals_s1_write -> pio_signals:write_n
	wire  [31:0] mm_interconnect_0_pio_signals_s1_readdata;                 // pio_signals:readdata -> mm_interconnect_0:pio_signals_s1_readdata
	wire  [31:0] mm_interconnect_0_lan_rst_s1_writedata;                    // mm_interconnect_0:LAN_RST_s1_writedata -> LAN_RST:writedata
	wire   [1:0] mm_interconnect_0_lan_rst_s1_address;                      // mm_interconnect_0:LAN_RST_s1_address -> LAN_RST:address
	wire         mm_interconnect_0_lan_rst_s1_chipselect;                   // mm_interconnect_0:LAN_RST_s1_chipselect -> LAN_RST:chipselect
	wire         mm_interconnect_0_lan_rst_s1_write;                        // mm_interconnect_0:LAN_RST_s1_write -> LAN_RST:write_n
	wire  [31:0] mm_interconnect_0_lan_rst_s1_readdata;                     // LAN_RST:readdata -> mm_interconnect_0:LAN_RST_s1_readdata
	wire         irq_mapper_receiver0_irq;                                  // epcs:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // LAN:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_d_irq_irq;                                             // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [LAN:reset_n, LAN_CS:reset_n, LAN_NINT:reset_n, LAN_RST:reset_n, cpu:reset_n, epcs:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, onchip_mem:reset, rst_translator:in_reset, sysid:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, epcs:reset_req, onchip_mem:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                         // cpu:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [data32:reset_n, data32_in:reset_n, mm_interconnect_0:pio_time_reset_reset_bridge_in_reset_reset, pio_addr:reset_n, pio_count2:reset_n, pio_count3:reset_n, pio_count4:reset_n, pio_count:reset_n, pio_rdata:reset_n, pio_signals:reset_n, pio_signals_0:reset_n, pio_time:reset_n, pio_wdata:reset_n]

	sopc_epcs epcs (
		.clk           (clk),                                                 //               clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                     //             reset.reset_n
		.reset_req     (rst_controller_reset_out_reset_req),                  //                  .reset_req
		.address       (mm_interconnect_0_epcs_epcs_control_port_address),    // epcs_control_port.address
		.chipselect    (mm_interconnect_0_epcs_epcs_control_port_chipselect), //                  .chipselect
		.dataavailable (),                                                    //                  .dataavailable
		.endofpacket   (),                                                    //                  .endofpacket
		.read_n        (~mm_interconnect_0_epcs_epcs_control_port_read),      //                  .read_n
		.readdata      (mm_interconnect_0_epcs_epcs_control_port_readdata),   //                  .readdata
		.readyfordata  (),                                                    //                  .readyfordata
		.write_n       (~mm_interconnect_0_epcs_epcs_control_port_write),     //                  .write_n
		.writedata     (mm_interconnect_0_epcs_epcs_control_port_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver0_irq),                            //               irq.irq
		.dclk          (dclk_from_the_epcs),                                  //          external.export
		.sce           (sce_from_the_epcs),                                   //                  .export
		.sdo           (sdo_from_the_epcs),                                   //                  .export
		.data0         (data0_to_the_epcs)                                    //                  .export
	);

	sopc_jtag_uart jtag_uart (
		.clk            (clk),                                                       //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	sopc_LAN lan (
		.clk           (clk),                                               //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_lan_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_lan_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_lan_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_lan_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_lan_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_lan_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver2_irq),                          //              irq.irq
		.MISO          (MISO_to_the_LAN),                                   //         external.export
		.MOSI          (MOSI_from_the_LAN),                                 //                 .export
		.SCLK          (SCLK_from_the_LAN),                                 //                 .export
		.SS_n          (SS_n_from_the_LAN)                                  //                 .export
	);

	sopc_LAN_CS lan_cs (
		.clk        (clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_lan_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lan_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lan_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lan_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lan_cs_s1_readdata),   //                    .readdata
		.out_port   (out_port_from_the_LAN_CS)                // external_connection.export
	);

	sopc_LAN_NINT lan_nint (
		.clk      (clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_lan_nint_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_lan_nint_s1_readdata), //                    .readdata
		.in_port  (in_port_to_the_LAN_NINT)                 // external_connection.export
	);

	sopc_LAN_CS lan_rst (
		.clk        (clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_lan_rst_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lan_rst_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lan_rst_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lan_rst_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lan_rst_s1_readdata),   //                    .readdata
		.out_port   (out_port_from_the_LAN_RST)                // external_connection.export
	);

	sopc_onchip_mem onchip_mem (
		.clk        (clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_onchip_mem_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_mem_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_mem_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_mem_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_mem_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_mem_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_mem_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)          //       .reset_req
	);

	sopc_cpu cpu (
		.clk                                   (clk),                                                 //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	sopc_sysid sysid (
		.clock    (clk),                                            //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	sopc_pio_time pio_time (
		.clk      (clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_pio_time_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_time_s1_readdata), //                    .readdata
		.in_port  (time_export)                             // external_connection.export
	);

	sopc_pio_time pio_count (
		.clk      (clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_pio_count_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_count_s1_readdata), //                    .readdata
		.in_port  (ch1_count_export)                         // external_connection.export
	);

	sopc_pio_addr pio_addr (
		.clk        (clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_pio_addr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_addr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_addr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_addr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_addr_s1_readdata),   //                    .readdata
		.out_port   (addr_export)                               // external_connection.export
	);

	sopc_pio_addr pio_wdata (
		.clk        (clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_wdata_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_wdata_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_wdata_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_wdata_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_wdata_s1_readdata),   //                    .readdata
		.out_port   (wdata_export)                               // external_connection.export
	);

	sopc_pio_rdata pio_rdata (
		.clk      (clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_pio_rdata_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_rdata_s1_readdata), //                    .readdata
		.in_port  (rdata_export)                             // external_connection.export
	);

	sopc_pio_addr pio_signals (
		.clk        (clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_signals_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_signals_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_signals_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_signals_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_signals_s1_readdata),   //                    .readdata
		.out_port   (signals_export)                               // external_connection.export
	);

	sopc_pio_rdata pio_signals_0 (
		.clk      (clk),                                         //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_pio_signals_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_signals_0_s1_readdata), //                    .readdata
		.in_port  (status_export)                                // external_connection.export
	);

	sopc_data32 data32 (
		.clk        (clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_data32_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_data32_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_data32_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_data32_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_data32_s1_readdata),   //                    .readdata
		.out_port   (wdata32_export)                          // external_connection.export
	);

	sopc_data32 data32_in (
		.clk        (clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_data32_in_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_data32_in_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_data32_in_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_data32_in_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_data32_in_s1_readdata),   //                    .readdata
		.out_port   (rdata32_export)                             // external_connection.export
	);

	sopc_pio_time pio_count2 (
		.clk      (clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_pio_count2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_count2_s1_readdata), //                    .readdata
		.in_port  (ch2_count_export)                          // external_connection.export
	);

	sopc_pio_time pio_count3 (
		.clk      (clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_pio_count3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_count3_s1_readdata), //                    .readdata
		.in_port  (ch3_count_export)                          // external_connection.export
	);

	sopc_pio_time pio_count4 (
		.clk      (clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_pio_count4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_count4_s1_readdata), //                    .readdata
		.in_port  (ch4_count_export)                          // external_connection.export
	);

	sopc_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                (clk),                                                       //                              clk_clk.clk
		.cpu_reset_n_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                            //    cpu_reset_n_reset_bridge_in_reset.reset
		.pio_time_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                        // pio_time_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                    (cpu_data_master_address),                                   //                      cpu_data_master.address
		.cpu_data_master_waitrequest                (cpu_data_master_waitrequest),                               //                                     .waitrequest
		.cpu_data_master_byteenable                 (cpu_data_master_byteenable),                                //                                     .byteenable
		.cpu_data_master_read                       (cpu_data_master_read),                                      //                                     .read
		.cpu_data_master_readdata                   (cpu_data_master_readdata),                                  //                                     .readdata
		.cpu_data_master_write                      (cpu_data_master_write),                                     //                                     .write
		.cpu_data_master_writedata                  (cpu_data_master_writedata),                                 //                                     .writedata
		.cpu_data_master_debugaccess                (cpu_data_master_debugaccess),                               //                                     .debugaccess
		.cpu_instruction_master_address             (cpu_instruction_master_address),                            //               cpu_instruction_master.address
		.cpu_instruction_master_waitrequest         (cpu_instruction_master_waitrequest),                        //                                     .waitrequest
		.cpu_instruction_master_read                (cpu_instruction_master_read),                               //                                     .read
		.cpu_instruction_master_readdata            (cpu_instruction_master_readdata),                           //                                     .readdata
		.cpu_jtag_debug_module_address              (mm_interconnect_0_cpu_jtag_debug_module_address),           //                cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                (mm_interconnect_0_cpu_jtag_debug_module_write),             //                                     .write
		.cpu_jtag_debug_module_read                 (mm_interconnect_0_cpu_jtag_debug_module_read),              //                                     .read
		.cpu_jtag_debug_module_readdata             (mm_interconnect_0_cpu_jtag_debug_module_readdata),          //                                     .readdata
		.cpu_jtag_debug_module_writedata            (mm_interconnect_0_cpu_jtag_debug_module_writedata),         //                                     .writedata
		.cpu_jtag_debug_module_byteenable           (mm_interconnect_0_cpu_jtag_debug_module_byteenable),        //                                     .byteenable
		.cpu_jtag_debug_module_waitrequest          (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),       //                                     .waitrequest
		.cpu_jtag_debug_module_debugaccess          (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),       //                                     .debugaccess
		.data32_s1_address                          (mm_interconnect_0_data32_s1_address),                       //                            data32_s1.address
		.data32_s1_write                            (mm_interconnect_0_data32_s1_write),                         //                                     .write
		.data32_s1_readdata                         (mm_interconnect_0_data32_s1_readdata),                      //                                     .readdata
		.data32_s1_writedata                        (mm_interconnect_0_data32_s1_writedata),                     //                                     .writedata
		.data32_s1_chipselect                       (mm_interconnect_0_data32_s1_chipselect),                    //                                     .chipselect
		.data32_in_s1_address                       (mm_interconnect_0_data32_in_s1_address),                    //                         data32_in_s1.address
		.data32_in_s1_write                         (mm_interconnect_0_data32_in_s1_write),                      //                                     .write
		.data32_in_s1_readdata                      (mm_interconnect_0_data32_in_s1_readdata),                   //                                     .readdata
		.data32_in_s1_writedata                     (mm_interconnect_0_data32_in_s1_writedata),                  //                                     .writedata
		.data32_in_s1_chipselect                    (mm_interconnect_0_data32_in_s1_chipselect),                 //                                     .chipselect
		.epcs_epcs_control_port_address             (mm_interconnect_0_epcs_epcs_control_port_address),          //               epcs_epcs_control_port.address
		.epcs_epcs_control_port_write               (mm_interconnect_0_epcs_epcs_control_port_write),            //                                     .write
		.epcs_epcs_control_port_read                (mm_interconnect_0_epcs_epcs_control_port_read),             //                                     .read
		.epcs_epcs_control_port_readdata            (mm_interconnect_0_epcs_epcs_control_port_readdata),         //                                     .readdata
		.epcs_epcs_control_port_writedata           (mm_interconnect_0_epcs_epcs_control_port_writedata),        //                                     .writedata
		.epcs_epcs_control_port_chipselect          (mm_interconnect_0_epcs_epcs_control_port_chipselect),       //                                     .chipselect
		.jtag_uart_avalon_jtag_slave_address        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //          jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                     .write
		.jtag_uart_avalon_jtag_slave_read           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                     .read
		.jtag_uart_avalon_jtag_slave_readdata       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                     .readdata
		.jtag_uart_avalon_jtag_slave_writedata      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                     .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                     .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                     .chipselect
		.LAN_spi_control_port_address               (mm_interconnect_0_lan_spi_control_port_address),            //                 LAN_spi_control_port.address
		.LAN_spi_control_port_write                 (mm_interconnect_0_lan_spi_control_port_write),              //                                     .write
		.LAN_spi_control_port_read                  (mm_interconnect_0_lan_spi_control_port_read),               //                                     .read
		.LAN_spi_control_port_readdata              (mm_interconnect_0_lan_spi_control_port_readdata),           //                                     .readdata
		.LAN_spi_control_port_writedata             (mm_interconnect_0_lan_spi_control_port_writedata),          //                                     .writedata
		.LAN_spi_control_port_chipselect            (mm_interconnect_0_lan_spi_control_port_chipselect),         //                                     .chipselect
		.LAN_CS_s1_address                          (mm_interconnect_0_lan_cs_s1_address),                       //                            LAN_CS_s1.address
		.LAN_CS_s1_write                            (mm_interconnect_0_lan_cs_s1_write),                         //                                     .write
		.LAN_CS_s1_readdata                         (mm_interconnect_0_lan_cs_s1_readdata),                      //                                     .readdata
		.LAN_CS_s1_writedata                        (mm_interconnect_0_lan_cs_s1_writedata),                     //                                     .writedata
		.LAN_CS_s1_chipselect                       (mm_interconnect_0_lan_cs_s1_chipselect),                    //                                     .chipselect
		.LAN_NINT_s1_address                        (mm_interconnect_0_lan_nint_s1_address),                     //                          LAN_NINT_s1.address
		.LAN_NINT_s1_readdata                       (mm_interconnect_0_lan_nint_s1_readdata),                    //                                     .readdata
		.LAN_RST_s1_address                         (mm_interconnect_0_lan_rst_s1_address),                      //                           LAN_RST_s1.address
		.LAN_RST_s1_write                           (mm_interconnect_0_lan_rst_s1_write),                        //                                     .write
		.LAN_RST_s1_readdata                        (mm_interconnect_0_lan_rst_s1_readdata),                     //                                     .readdata
		.LAN_RST_s1_writedata                       (mm_interconnect_0_lan_rst_s1_writedata),                    //                                     .writedata
		.LAN_RST_s1_chipselect                      (mm_interconnect_0_lan_rst_s1_chipselect),                   //                                     .chipselect
		.onchip_mem_s1_address                      (mm_interconnect_0_onchip_mem_s1_address),                   //                        onchip_mem_s1.address
		.onchip_mem_s1_write                        (mm_interconnect_0_onchip_mem_s1_write),                     //                                     .write
		.onchip_mem_s1_readdata                     (mm_interconnect_0_onchip_mem_s1_readdata),                  //                                     .readdata
		.onchip_mem_s1_writedata                    (mm_interconnect_0_onchip_mem_s1_writedata),                 //                                     .writedata
		.onchip_mem_s1_byteenable                   (mm_interconnect_0_onchip_mem_s1_byteenable),                //                                     .byteenable
		.onchip_mem_s1_chipselect                   (mm_interconnect_0_onchip_mem_s1_chipselect),                //                                     .chipselect
		.onchip_mem_s1_clken                        (mm_interconnect_0_onchip_mem_s1_clken),                     //                                     .clken
		.pio_addr_s1_address                        (mm_interconnect_0_pio_addr_s1_address),                     //                          pio_addr_s1.address
		.pio_addr_s1_write                          (mm_interconnect_0_pio_addr_s1_write),                       //                                     .write
		.pio_addr_s1_readdata                       (mm_interconnect_0_pio_addr_s1_readdata),                    //                                     .readdata
		.pio_addr_s1_writedata                      (mm_interconnect_0_pio_addr_s1_writedata),                   //                                     .writedata
		.pio_addr_s1_chipselect                     (mm_interconnect_0_pio_addr_s1_chipselect),                  //                                     .chipselect
		.pio_count_s1_address                       (mm_interconnect_0_pio_count_s1_address),                    //                         pio_count_s1.address
		.pio_count_s1_readdata                      (mm_interconnect_0_pio_count_s1_readdata),                   //                                     .readdata
		.pio_count2_s1_address                      (mm_interconnect_0_pio_count2_s1_address),                   //                        pio_count2_s1.address
		.pio_count2_s1_readdata                     (mm_interconnect_0_pio_count2_s1_readdata),                  //                                     .readdata
		.pio_count3_s1_address                      (mm_interconnect_0_pio_count3_s1_address),                   //                        pio_count3_s1.address
		.pio_count3_s1_readdata                     (mm_interconnect_0_pio_count3_s1_readdata),                  //                                     .readdata
		.pio_count4_s1_address                      (mm_interconnect_0_pio_count4_s1_address),                   //                        pio_count4_s1.address
		.pio_count4_s1_readdata                     (mm_interconnect_0_pio_count4_s1_readdata),                  //                                     .readdata
		.pio_rdata_s1_address                       (mm_interconnect_0_pio_rdata_s1_address),                    //                         pio_rdata_s1.address
		.pio_rdata_s1_readdata                      (mm_interconnect_0_pio_rdata_s1_readdata),                   //                                     .readdata
		.pio_signals_s1_address                     (mm_interconnect_0_pio_signals_s1_address),                  //                       pio_signals_s1.address
		.pio_signals_s1_write                       (mm_interconnect_0_pio_signals_s1_write),                    //                                     .write
		.pio_signals_s1_readdata                    (mm_interconnect_0_pio_signals_s1_readdata),                 //                                     .readdata
		.pio_signals_s1_writedata                   (mm_interconnect_0_pio_signals_s1_writedata),                //                                     .writedata
		.pio_signals_s1_chipselect                  (mm_interconnect_0_pio_signals_s1_chipselect),               //                                     .chipselect
		.pio_signals_0_s1_address                   (mm_interconnect_0_pio_signals_0_s1_address),                //                     pio_signals_0_s1.address
		.pio_signals_0_s1_readdata                  (mm_interconnect_0_pio_signals_0_s1_readdata),               //                                     .readdata
		.pio_time_s1_address                        (mm_interconnect_0_pio_time_s1_address),                     //                          pio_time_s1.address
		.pio_time_s1_readdata                       (mm_interconnect_0_pio_time_s1_readdata),                    //                                     .readdata
		.pio_wdata_s1_address                       (mm_interconnect_0_pio_wdata_s1_address),                    //                         pio_wdata_s1.address
		.pio_wdata_s1_write                         (mm_interconnect_0_pio_wdata_s1_write),                      //                                     .write
		.pio_wdata_s1_readdata                      (mm_interconnect_0_pio_wdata_s1_readdata),                   //                                     .readdata
		.pio_wdata_s1_writedata                     (mm_interconnect_0_pio_wdata_s1_writedata),                  //                                     .writedata
		.pio_wdata_s1_chipselect                    (mm_interconnect_0_pio_wdata_s1_chipselect),                 //                                     .chipselect
		.sysid_control_slave_address                (mm_interconnect_0_sysid_control_slave_address),             //                  sysid_control_slave.address
		.sysid_control_slave_readdata               (mm_interconnect_0_sysid_control_slave_readdata)             //                                     .readdata
	);

	sopc_irq_mapper irq_mapper (
		.clk           (clk),                            //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.clk            (clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
